
// データ幅は16bit
`define DATA_WIDTH 16

// データパス
`define DataPath logic [ `DATA_WIDTH-1:0 ]
